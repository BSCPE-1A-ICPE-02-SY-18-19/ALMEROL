CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 5 110 10
176 80 1278 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 846 4 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
43530.3 0
0
6 74LS48
188 793 151 0 14 29
0 4 7 6 5 18 19 10 11 12
13 14 15 16 20
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
391 0 0
2
43530.3 0
0
9 CC 7-Seg~
183 846 58 0 17 19
10 16 15 14 13 12 11 10 21 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3124 0 0
2
43530.3 1
0
9 2-In AND~
219 622 112 0 3 22
0 9 7 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3421 0 0
2
43530.3 2
0
9 2-In AND~
219 484 111 0 3 22
0 5 6 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8157 0 0
2
43530.3 3
0
2 +V
167 258 167 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
43530.3 4
0
7 Pulser~
4 858 434 0 10 12
0 22 3 23 3 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
5.89883e-315 0
0
6 74112~
219 681 276 0 7 32
0 8 17 3 17 8 24 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
7361 0 0
2
5.89883e-315 5.26354e-315
0
6 74112~
219 542 276 0 7 32
0 8 9 3 9 8 25 7
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4747 0 0
2
5.89883e-315 5.30499e-315
0
6 74112~
219 394 278 0 7 32
0 8 5 3 5 8 26 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
972 0 0
2
5.89883e-315 5.32571e-315
0
6 74112~
219 261 277 0 7 32
0 8 27 3 28 8 29 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3472 0 0
2
5.89883e-315 5.34643e-315
0
37
2 0 3 0 0 4096 0 7 0 0 37 4
828 434
828 349
824 349
824 364
1 9 2 0 0 4224 0 1 3 0 0 4
846 12
846 24
846 24
846 16
7 1 4 0 0 8320 0 8 2 0 0 4
705 240
753 240
753 115
761 115
0 4 5 0 0 8320 0 0 2 27 0 3
330 241
330 142
761 142
0 3 6 0 0 12416 0 0 2 34 0 4
439 240
458 240
458 133
761 133
0 2 7 0 0 12416 0 0 2 33 0 4
590 241
621 241
621 124
761 124
0 0 8 0 0 4096 0 0 0 10 24 2
633 289
633 189
0 0 8 0 0 0 0 0 0 11 24 2
469 289
469 189
0 0 8 0 0 0 0 0 0 24 12 2
312 189
312 289
5 5 8 0 0 0 0 9 8 0 0 6
542 288
633 288
633 289
633 289
633 288
681 288
5 5 8 0 0 0 0 10 9 0 0 4
394 290
469 290
469 288
542 288
5 5 8 0 0 0 0 11 10 0 0 4
261 289
312 289
312 290
394 290
2 0 9 0 0 12288 0 9 0 0 14 4
518 240
515 240
515 241
505 241
4 3 9 0 0 8320 0 9 5 0 0 3
518 258
505 258
505 111
7 7 10 0 0 4224 0 2 3 0 0 3
825 115
861 115
861 94
8 6 11 0 0 4224 0 2 3 0 0 3
825 124
855 124
855 94
9 5 12 0 0 8320 0 2 3 0 0 3
825 133
849 133
849 94
10 4 13 0 0 8320 0 2 3 0 0 3
825 142
843 142
843 94
11 3 14 0 0 8320 0 2 3 0 0 3
825 151
837 151
837 94
12 2 15 0 0 8320 0 2 3 0 0 3
825 160
831 160
831 94
13 1 16 0 0 4224 0 2 3 0 0 2
825 169
825 94
1 0 8 0 0 0 0 9 0 0 24 4
542 213
542 201
549 201
549 189
1 0 8 0 0 0 0 10 0 0 24 4
394 215
394 196
392 196
392 189
1 0 8 0 0 8320 0 8 0 0 25 3
681 213
681 189
258 189
1 1 8 0 0 0 0 11 6 0 0 4
261 214
261 189
258 189
258 176
2 0 5 0 0 0 0 10 0 0 27 4
370 242
361 242
361 241
355 241
7 0 5 0 0 0 0 11 0 0 28 2
285 241
355 241
1 4 5 0 0 0 0 5 10 0 0 4
460 102
355 102
355 260
370 260
3 0 3 0 0 0 0 11 0 0 37 3
231 250
206 250
206 321
3 1 9 0 0 0 0 5 4 0 0 3
505 111
505 103
598 103
2 0 17 0 0 12288 0 8 0 0 32 4
657 240
663 240
663 241
653 241
3 4 17 0 0 8320 0 4 8 0 0 4
643 112
653 112
653 258
657 258
7 2 7 0 0 0 0 9 4 0 0 6
566 240
590 240
590 241
590 241
590 121
598 121
2 7 6 0 0 0 0 5 10 0 0 4
460 120
439 120
439 242
418 242
3 0 3 0 0 0 0 9 0 0 37 3
512 249
487 249
487 321
3 0 3 0 0 0 0 10 0 0 37 3
364 251
340 251
340 321
4 3 3 0 0 8336 0 7 8 0 0 7
888 434
888 364
206 364
206 321
641 321
641 249
651 249
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
